library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ControlUnit is
port (CLK: in std_logic;
		Word: in std_logic_vector(15 downto 0);
		NZCV: in std_lOGIC_vector(3 downto 0);
		
		FLAGS: out std_logic;
		 SEL: out STD_LOGIC_vector(4 downto 0);--ALU
		 WE: out std_logic;--banco de registros
		 RE: out std_logic;--banco de registros
		 RdAdd: out std_logic_vector(3 downto 0);
		 RnAdd: out std_logic_vector(3 downto 0);--banco de registros
		 RmAdd: out std_logic_vector(3 downto 0);--banco de registros
		 WR: out std_logic; --RAM
		 
		 MUX_SEL: out std_logic;
		 read_rom: out std_logic;
		 ARLOAD: OUT STD_LOGIC;
		 ZLOAD_1: OUT STD_LOGIC;
		 ZLOAD_2: OUT STD_LOGIC;
		 ZLOAD_3: OUT STD_LOGIC;
		 IMM: OUT STD_LOGIC_vector(31 DOWNTO 0);
		 PCINC: OUT STD_LOGIC;
		 CarryEn: out std_logic
		 
		);
end ControlUnit;
	
architecture RTL of ControlUnit is
signal IR: std_logic_vector(15 downto 0);
signal IRload: std_logic;

signal IR2: std_logic_vector(15 downto 0);
signal IRload2: std_logic;

signal BIFURCATION: std_lOGIC_vector(3 downto 0);


--SENALES DE CONTROL--
signal estados: std_logic_vector(127 downto 0);
SIGNAL COUNTER: STD_LOGIC_VECTOR(6 DOWNTO 0);
signal CTRLINC: STD_LOGIC;
SIGNAL CTRLCLEAR: STD_LOGIC;
signal CTRLOAD: STD_LOGIC;


signal FETCH1,FETCH2,FETCH3: STD_LOGIC;
signal ALU1,ALU2: STD_LOGIC;
signal STR1,STR2,STR3,STR4,STR5: STD_LOGIC;
SIGNAL LOAD1,LOAD2,LOAD3,LOAD3T,LOAD4,LOAD5: STD_LOGIC;
signal MUL1,MUL2,MUL3,MUL4,MUL5,MUL6,MUL7,MUL8,MUL9,MUL10,MUL11,MUL12,MUL13,MUL14,MUL15,MUL16,MUL17,MUL18: STD_LOGIC;
signal BLX1,BLX2,BLX3,BLX4: STD_LOGIC;
signal BL1,BL2,BL3,BL4,BL5: STD_LOGIC;
signal PUSH1,PUSH2,PUSH3,PUSH4,PUSH5,PUSH6,PUSH7,PUSH8,PUSH9,PUSH10,PUSH11,PUSH12,PUSH13,PUSH14,PUSH15:STD_LOGIC;
signal PUSH16,PUSH17,PUSH18,PUSH19,PUSH20,PUSH21,PUSH22,PUSH23,PUSH24,PUSH25,PUSH26,PUSH27,PUSH28,PUSH29,PUSH30:STD_LOGIC;
signal PUSH31,PUSH32,PUSH33,PUSH34,PUSH35,PUSH36,PUSH37,PUSH38,PUSH39,PUSH40,PUSH41,PUSH42,PUSH43,PUSH44,PUSH45:STD_LOGIC;
signal POP1,POP2,POP3,POP4,POP5,POP6,POP7,POP8,POP9,POP10,POP11,POP12,POP13,POP14,POP15:STD_LOGIC;
signal POP16,POP17,POP18,POP19,POP20,POP21,POP22,POP23,POP24,POP25,POP26,POP27,POP28,POP29,POP30:STD_LOGIC;
signal POP31,POP32,POP33,POP34,POP35,POP36,POP37,POP38:STD_LOGIC;

begin

CONTROLLER: PROCESS(CLK) BEGin
if clk'event and clk='0' then

	IF CTRLINC='1' THEN--COUNTER; SALIDA DEL CONTADOR PARA PROVEER AL DECODIFICADOR
			COUNTER<=COUNTER+'1';
	ELSIF CTRLCLEAR='1' THEN
			COUNTER<=(OTHERS=>'0');
	ELSIF CTRLOAD='1' THEN
			IF (BIFURCATION="0000" OR BIFURCATION="0001") THEN
				COUNTER<="0000011";
			ELSIF BIFURCATION="0010" THEN
				COUNTER<="0010000";
			ELSIF BIFURCATION="0011" THEN
				COUNTER<="0000101";
			ELSIF (BIFURCATION="0100" OR BIFURCATION="0101") THEN
				COUNTER<="0001010";
			ELSIF (BIFURCATION="0110") THEN
				COUNTER<="0100010";
			ELSIF (BIFURCATION="0111") THEN
				COUNTER<="0100110";
			ELSIF (BIFURCATION="1000") THEN
				IF(FETCH3='1')THEN
					COUNTER<="0101011";
				ELSIF(PUSH1='1')THEN
					COUNTER<="0110000";
				ELSIF(PUSH6='1')THEN
					COUNTER<="0110101";
				ELSIF(PUSH11='1')THEN
					COUNTER<="0111010";
				ELSIF(PUSH16='1')THEN
					COUNTER<="0111111";
				ELSIF(PUSH21='1')THEN
					COUNTER<="1000100";
				ELSIF(PUSH26='1')THEN
					COUNTER<="1001001";
				ELSIF(PUSH31='1')THEN
					COUNTER<="1001110";
				ELSIF(PUSH36='1')THEN
					COUNTER<="1010011";
				ELSE
					COUNTER<="0000000";
				END IF;
			ELSIF (BIFURCATION="1001") THEN
				IF(FETCH3='1')THEN
					COUNTER<="1011000";
				ELSIF(POP3='1')THEN
					COUNTER<="1011110";
				ELSIF(POP7='1')THEN
					COUNTER<="1100010";
				ELSIF(POP11='1')THEN
					COUNTER<="1100110";
				ELSIF(POP15='1')THEN
					COUNTER<="1101010";
				ELSIF(POP19='1')THEN
					COUNTER<="1101110";
				ELSIF(POP23='1')THEN
					COUNTER<="1110010";
				ELSIF(POP27='1')THEN
					COUNTER<="1110110";
				ELSIF(POP31='1')THEN
					COUNTER<="1111010";
				ELSE
					COUNTER<="0000000";
				END IF;
			ELSE
				COUNTER<="0000000";
			END IF;
	END IF;
	
else null;
end if;
end process;


ESTADOS<="00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001" when COUNTER="0000000" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010" WHEN COUNTER="0000001" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100" WHEN COUNTER="0000010" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000" WHEN COUNTER="0000011" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000" when COUNTER="0000100" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000" WHEN COUNTER="0000101" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000" WHEN COUNTER="0000110" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000" WHEN COUNTER="0000111" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000" when COUNTER="0001000" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000" WHEN COUNTER="0001001" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000" WHEN COUNTER="0001010" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000" WHEN COUNTER="0001011" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000" when COUNTER="0001100" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000" WHEN COUNTER="0001101" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000" WHEN COUNTER="0001110" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000" WHEN COUNTER="0001111" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000" when COUNTER="0010000" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000" WHEN COUNTER="0010001" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000" WHEN COUNTER="0010010" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000" WHEN COUNTER="0010011" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000" when COUNTER="0010100" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000" WHEN COUNTER="0010101" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000" WHEN COUNTER="0010110" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000" WHEN COUNTER="0010111" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000" when COUNTER="0011000" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000" WHEN COUNTER="0011001" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000" WHEN COUNTER="0011010" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000" WHEN COUNTER="0011011" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000" when COUNTER="0011100" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000" WHEN COUNTER="0011101" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000" WHEN COUNTER="0011110" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000" WHEN COUNTER="0011111" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000" when COUNTER="0100000" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000" WHEN COUNTER="0100001" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000" WHEN COUNTER="0100010" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000" WHEN COUNTER="0100011" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000" when COUNTER="0100100" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000" WHEN COUNTER="0100101" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000" WHEN COUNTER="0100110" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000" WHEN COUNTER="0100111" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000" when COUNTER="0101000" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000" WHEN COUNTER="0101001" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000" WHEN COUNTER="0101010" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000" WHEN COUNTER="0101011" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000" when COUNTER="0101100" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000" WHEN COUNTER="0101101" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000" WHEN COUNTER="0101110" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000" WHEN COUNTER="0101111" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000" when COUNTER="0110000" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000" WHEN COUNTER="0110001" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000" WHEN COUNTER="0110010" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000" WHEN COUNTER="0110011" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000" when COUNTER="0110100" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000" WHEN COUNTER="0110101" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000" WHEN COUNTER="0110110" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000" WHEN COUNTER="0110111" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000" when COUNTER="0111000" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="0111001" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="0111010" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="0111011" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000" when COUNTER="0111100" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="0111101" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="0111110" ELSE
			"00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="0111111" ELSE
			"00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000" when COUNTER="1000000" ELSE
			"00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1000001" ELSE
			"00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1000010" ELSE
			"00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1000011" ELSE
			"00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000" when COUNTER="1000100" ELSE
			"00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1000101" ELSE
			"00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1000110" ELSE
			"00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1000111" ELSE
			"00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000" when COUNTER="1001000" ELSE
			"00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1001001" ELSE
			"00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1001010" ELSE
			"00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1001011" ELSE
			"00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000" when COUNTER="1001100" ELSE
			"00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1001101" ELSE
			"00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1001110" ELSE
			"00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1001111" ELSE
			"00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000" when COUNTER="1010000" ELSE
			"00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1010001" ELSE
			"00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1010010" ELSE
			"00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1010011" ELSE
			"00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000" when COUNTER="1010100" ELSE
			"00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1010101" ELSE
			"00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1010110" ELSE
			"00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1010111" ELSE
			"00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" when COUNTER="1011000" ELSE
			"00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1011001" ELSE
			"00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1011010" ELSE
			"00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1011011" ELSE
			"00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" when COUNTER="1011100" ELSE
			"00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1011101" ELSE
			"00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1011110" ELSE
			"00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1011111" ELSE
			"00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" when COUNTER="1100000" ELSE
			"00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1100001" ELSE
			"00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1100010" ELSE
			"00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1100011" ELSE
			"00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" when COUNTER="1100100" ELSE
			"00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1100101" ELSE
			"00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1100110" ELSE
			"00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1100111" ELSE
			"00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" when COUNTER="1101000" ELSE
			"00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1101001" ELSE
			"00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1101010" ELSE
			"00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1101011" ELSE
			"00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" when COUNTER="1101100" ELSE
			"00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1101101" ELSE
			"00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1101110" ELSE
			"00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1101111" ELSE
			"00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" when COUNTER="1110000" ELSE
			"00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1110001" ELSE
			"00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1110010" ELSE
			"00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1110011" ELSE
			"00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" when COUNTER="1110100" ELSE
			"00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1110101" ELSE
			"00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1110110" ELSE
			"00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1110111" ELSE
			"00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" when COUNTER="1111000" ELSE
			"00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1111001" ELSE
			"00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1111010" ELSE
			"00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1111011" ELSE
			"00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" when COUNTER="1111100" ELSE
			"00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1111101" ELSE
			"01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1111110" ELSE
			"10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" WHEN COUNTER="1111111" ELSE
			"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

FETCH1<=ESTADOS(0);
FETCH2<=ESTADOS(1);
FETCH3<=ESTADOS(2);

ALU1<=ESTADOS(3);
ALU2<=ESTADOS(4);

STR1<=ESTADOS(5);
STR2<=ESTADOS(6);
STR3<=ESTADOS(7);
STR4<=ESTADOS(8);
STR5<=ESTADOS(9);

LOAD1<=ESTADOS(10);
LOAD2<=ESTADOS(11);
LOAD3<=ESTADOS(12);
LOAD3T<=ESTADOS(13);
LOAD4<=ESTADOS(14);
LOAD5<=ESTADOS(15);

MUL1<=ESTADOS(16);
MUL2<=ESTADOS(17);
MUL3<=ESTADOS(18);
MUL4<=ESTADOS(19);
MUL5<=ESTADOS(20);
MUL6<=ESTADOS(21);
MUL7<=ESTADOS(22);
MUL8<=ESTADOS(23);
MUL9<=ESTADOS(24);
MUL10<=ESTADOS(25);
MUL11<=ESTADOS(26);
MUL12<=ESTADOS(27);
MUL13<=ESTADOS(28);
MUL14<=ESTADOS(29);
MUL15<=ESTADOS(30);
MUL16<=ESTADOS(31);
MUL17<=ESTADOS(32);
MUL18<=ESTADOS(33);

BLX1<=ESTADOS(34);
BLX2<=ESTADOS(35);
BLX3<=ESTADOS(36);
BLX4<=ESTADOS(37);

BL1<=ESTADOS(38);
BL2<=ESTADOS(39);
BL3<=ESTADOS(40);
BL4<=ESTADOS(41);
BL5<=ESTADOS(42);

PUSH1<=ESTADOS(43);
PUSH2<=ESTADOS(44);
PUSH3<=ESTADOS(45);
PUSH4<=ESTADOS(46);
PUSH5<=ESTADOS(47);
PUSH6<=ESTADOS(48);
PUSH7<=ESTADOS(49);
PUSH8<=ESTADOS(50);
PUSH9<=ESTADOS(51);
PUSH10<=ESTADOS(52);
PUSH11<=ESTADOS(53);
PUSH12<=ESTADOS(54);
PUSH13<=ESTADOS(55);
PUSH14<=ESTADOS(56);
PUSH15<=ESTADOS(57);
PUSH16<=ESTADOS(58);
PUSH17<=ESTADOS(59);
PUSH18<=ESTADOS(60);
PUSH19<=ESTADOS(61);
PUSH20<=ESTADOS(62);
PUSH21<=ESTADOS(63);
PUSH22<=ESTADOS(64);
PUSH23<=ESTADOS(65);
PUSH24<=ESTADOS(66);
PUSH25<=ESTADOS(67);
PUSH26<=ESTADOS(68);
PUSH27<=ESTADOS(69);
PUSH28<=ESTADOS(70);
PUSH29<=ESTADOS(71);
PUSH30<=ESTADOS(72);
PUSH31<=ESTADOS(73);
PUSH32<=ESTADOS(74);
PUSH33<=ESTADOS(75);
PUSH34<=ESTADOS(76);
PUSH35<=ESTADOS(77);
PUSH36<=ESTADOS(78);
PUSH37<=ESTADOS(79);
PUSH38<=ESTADOS(80);
PUSH39<=ESTADOS(81);
PUSH40<=ESTADOS(82);
PUSH41<=ESTADOS(83);
PUSH42<=ESTADOS(84);
PUSH43<=ESTADOS(85);
PUSH44<=ESTADOS(86);
PUSH45<=ESTADOS(87);

POP1<=ESTADOS(88);
POP2<=ESTADOS(89);
POP3<=ESTADOS(90);
POP4<=ESTADOS(91);
POP5<=ESTADOS(92);
POP6<=ESTADOS(93);
POP7<=ESTADOS(94);
POP8<=ESTADOS(95);
POP9<=ESTADOS(96);
POP10<=ESTADOS(97);
POP11<=ESTADOS(98);
POP12<=ESTADOS(99);
POP13<=ESTADOS(100);
POP14<=ESTADOS(101);
POP15<=ESTADOS(102);
POP16<=ESTADOS(103);
POP17<=ESTADOS(104);
POP18<=ESTADOS(105);
POP19<=ESTADOS(106);
POP20<=ESTADOS(107);
POP21<=ESTADOS(108);
POP22<=ESTADOS(109);
POP23<=ESTADOS(110);
POP24<=ESTADOS(111);
POP25<=ESTADOS(112);
POP26<=ESTADOS(113);
POP27<=ESTADOS(114);
POP28<=ESTADOS(115);
POP29<=ESTADOS(116);
POP30<=ESTADOS(117);
POP31<=ESTADOS(118);
POP32<=ESTADOS(119);
POP33<=ESTADOS(120);
POP34<=ESTADOS(121);
POP35<=ESTADOS(122);
POP36<=ESTADOS(123);
POP37<=ESTADOS(124);
POP38<=ESTADOS(125);


ARLOAD<=FETCH1 OR BL1;
read_rom<=FETCH2 OR BL2;
PCINC<=FETCH2 OR BL2;
IRLOAD<=FETCH3;
IRLOAD2<=BL3;

RE<=ALU1 OR STR1 OR STR3 OR LOAD1 OR LOAD4 OR MUL1 OR BLX1 OR BLX3 OR BL1 OR BL4 OR PUSH1 OR PUSH3 OR PUSH6 OR PUSH8 OR PUSH11 OR PUSH13 OR PUSH16 OR PUSH18 OR PUSH21 OR PUSH23 OR PUSH26 OR PUSH28 OR PUSH31 OR PUSH33 OR PUSH36 OR PUSH38 OR PUSH41 OR PUSH43 OR POP1 OR POP3 OR POP7 OR POP11 OR POP15 OR POP19 OR POP23 OR POP27 OR POP31 OR POP35;
ZLOAD_1<=ALU2 OR STR2 OR STR4 OR STR5 OR LOAD2 OR LOAD5 OR MUL18 OR BLX2 OR BLX4 OR BL2 OR BL5 OR PUSH4 OR PUSH5 OR PUSH9 OR PUSH10 OR PUSH14 OR PUSH15 OR PUSH19 OR PUSH20 OR PUSH24 OR PUSH25 OR PUSH29 OR PUSH30 OR PUSH34 OR PUSH35 OR PUSH39 OR PUSH40 OR PUSH44 OR PUSH45 OR PUSH2 OR PUSH7 OR PUSH12 OR PUSH17 OR PUSH22 OR PUSH27 OR PUSH32 OR PUSH37 OR PUSH42 OR POP2 OR POP4 OR POP8 OR POP12 OR POP16 OR POP20 OR POP24 OR POP28 OR POP32 OR POP36 ;
ZLOAD_2<=STR2 OR LOAD2 OR PUSH2 OR PUSH7 OR PUSH12 OR PUSH17 OR PUSH22 OR PUSH27 OR PUSH32 OR PUSH37 OR PUSH42 OR POP4 OR POP8 OR POP12 OR POP16 OR POP20 OR POP24 OR POP28 OR POP32 OR POP36 ;
ZLOAD_3<=STR5 OR LOAD3 OR LOAD3T OR STR4 OR PUSH4 OR PUSH5 OR PUSH9 OR PUSH10 OR PUSH14 OR PUSH15 OR PUSH19 OR PUSH20 OR PUSH24 OR PUSH25 OR PUSH29 OR PUSH30 OR PUSH34 OR PUSH35 OR PUSH39 OR PUSH40 OR PUSH44 OR PUSH45 OR POP6 OR POP10 OR POP14 OR POP18 OR POP22 OR POP26 OR POP30 OR POP34 OR POP38 OR POP5 OR POP9 OR POP13 OR POP17 OR POP21 OR POP25 OR POP29 OR POP33 OR POP37;

WE<=ALU2 OR LOAD3T OR LOAD5 OR MUL18 OR BLX2 OR BLX4 OR BL2 OR BL5 OR PUSH2 OR PUSH7 OR PUSH12 OR PUSH17 OR PUSH22 OR PUSH27 OR PUSH32 OR PUSH37 OR PUSH42 OR POP2 OR POP4 OR POP8 OR POP12 OR POP16 OR POP20 OR POP24 OR POP28 OR POP32 OR POP36 OR POP6 OR POP10 OR POP14 OR POP18 OR POP22 OR POP26 OR POP30 OR POP34 OR POP38;
WR<=STR4 OR STR5 OR PUSH4 OR PUSH5 OR PUSH9 OR PUSH10 OR PUSH14 OR PUSH15 OR PUSH19 OR PUSH20 OR PUSH24 OR PUSH25 OR PUSH29 OR PUSH30 OR PUSH34 OR PUSH35 OR PUSH39 OR PUSH40 OR PUSH44 OR PUSH45;

CTRLINC<=FETCH1 OR FETCH2 OR (ALU1 AND NOT(BIFURCATION(0))) OR STR1 OR STR2 OR STR3 OR STR4 OR LOAD1 OR LOAD2 OR LOAD3 OR (LOAD3T AND BIFURCATION(0)) OR LOAD4 OR MUL1 OR MUL2 OR MUL3 OR MUL4 OR MUL5 OR MUL6 OR MUL7 OR MUL8 OR MUL9 OR MUL10 OR MUL11 OR MUL12 OR MUL13 OR MUL14 OR MUL15 OR MUL16 OR MUL17 OR BLX1 OR BLX2 OR BLX3 OR BL1 OR BL2 OR BL3 OR BL4 OR (PUSH1 AND IR(0)) OR PUSH2 OR PUSH3 OR PUSH4 OR PUSH5 OR (PUSH6 AND IR(1)) OR PUSH7 OR PUSH8 OR PUSH9 OR PUSH10 OR(PUSH11 AND IR(2)) OR PUSH12 OR PUSH13 OR PUSH14 OR PUSH15 OR (PUSH16 AND IR(3)) OR PUSH17 OR PUSH18 OR PUSH19 OR PUSH20 OR (PUSH21 AND IR(4)) OR PUSH22 OR PUSH23 OR PUSH24 OR PUSH25 OR (PUSH26 AND IR(5)) OR PUSH27 OR PUSH28 OR PUSH29 OR PUSH30 OR (PUSH31 AND IR(6)) OR PUSH32 OR PUSH33 OR PUSH34 OR PUSH35 OR (PUSH36 AND IR(7)) OR PUSH37 OR PUSH38 OR PUSH39 OR PUSH40 OR (PUSH41 AND IR(8)) OR PUSH42 OR PUSH43 OR PUSH44 OR POP1 OR POP2 OR (POP3 AND IR(0)) OR POP4 OR POP5 OR POP6 OR (POP7 AND IR(1)) OR POP8 OR POP9 OR POP10 OR (POP11 AND IR(2)) OR POP12 OR POP13 OR POP14 OR (POP15 AND IR(3)) OR POP16 OR POP17 OR POP18 OR (POP19 AND IR(4)) OR POP20 OR POP21 OR POP22 OR (POP23 AND IR(5)) OR POP24 OR POP25 OR POP26 OR (POP27 AND IR(6)) OR POP28 OR POP29 OR POP30 OR (POP31 AND IR(7)) OR POP32 OR POP33 OR POP34 OR (POP35 AND IR(8)) OR POP36 OR POP37 ;
CTRLCLEAR<=ALU2 OR (ALU1 AND BIFURCATION(0)) OR STR5 OR LOAD5 OR (LOAD3T AND NOT(BIFURCATION(0))) OR MUL18 OR BLX4 OR BL5 OR PUSH45 OR (PUSH41 AND NOT(IR(8))) OR POP38 OR(POP35 AND NOT(IR(8)));
CTRLOAD<=FETCH3 OR (PUSH1 AND NOT(IR(0))) OR (PUSH6 AND NOT(IR(1))) OR (PUSH11 AND NOT(IR(2))) OR (PUSH16 AND NOT(IR(3))) OR (PUSH21 AND NOT(IR(4))) OR (PUSH26 AND NOT(IR(5))) OR (PUSH31 AND NOT(IR(6))) OR (PUSH36 AND NOT(IR(7))) OR(POP3 AND NOT(IR(0))) OR(POP7 AND NOT(IR(1))) OR(POP11 AND NOT(IR(2))) OR(POP15 AND NOT(IR(3))) OR(POP19 AND NOT(IR(4))) OR(POP23 AND NOT(IR(5))) OR(POP27 AND NOT(IR(6))) OR(POP31 AND NOT(IR(7)));


process (clk) begin
if clk'event and clk='1' theN
	if IRLOAD='1' then
		IR<=word;
	else
		IR<=IR;
	end if;
else null;
end if;
end process;

process (clk) begin
if clk'event and clk='1' theN
	if IRLOAD2='1' then
		IR2<=word;
	else
		IR2<=IR2;
	end if;
else null;
end if;
end process;


---*****RECODIFICACION*****---
PROCESS(IR,ESTADOS) BEGin

	case IR(15 DOWNTO 14) is
		when "00" =>--Shift(immediate),add,subtract,move and compare
							 case IR(13 DOWNTO 11) is
									when "000" => SEL<="00110";--LSL(IMMEDIATE)
														 IMM<="000000000000000000000000000"&IR(10 DOWNTO 6);
														 MUX_SEL<='1';
														 Rmadd<='0'&IR(5 DOWNTO 3);
														 Rnadd<='0'&IR(5 DOWNTO 3);
														 Rdadd<='0'&IR(2 DOWNTO 0);
														 FLAGS<='1';
														 CarryEn<='1';
														 BIFURCATION<="0000";
														 
									when "001" => SEL<="00111";--LSR(IMMEDIATE)
														 IMM<="000000000000000000000000000"&IR(10 DOWNTO 6);
														 MUX_SEL<='1';
														 Rmadd<='0'&IR(5 DOWNTO 3);
														 Rnadd<='0'&IR(5 DOWNTO 3);
														 Rdadd<='0'&IR(2 DOWNTO 0);
														 FLAGS<='1';
														 CarryEn<='1';
														 BIFURCATION<="0000";
														 
									when "010" => SEL<="10000";--ASR(immEDIATE)
														 IMM<="000000000000000000000000000"&IR(10 DOWNTO 6);
														 MUX_SEL<='1';
														 Rmadd<='0'&IR(5 DOWNTO 3);
														 Rnadd<='0'&IR(5 DOWNTO 3);
														 Rdadd<='0'&IR(2 DOWNTO 0);
														 FLAGS<='1';
														 CarryEn<='1';
														 BIFURCATION<="0000";
									WHEN "011" =>
												CASE IR(13 DOWNTO 9) IS
													when "01100" => SEL<="00100";--ADD(register)T1
																		 MUX_SEL<='0';
																		 Rmadd<='0'&IR(8 DOWNTO 6);
																		 Rnadd<='0'&IR(5 DOWNTO 3);
																		 Rdadd<='0'&IR(2 DOWNTO 0);
																		 FLAGS<='1';
																		 CarryEn<='0';
																		 BIFURCATION<="0000";
																		 
													when "01101" => SEL<="00101";--SUB(register)
																		 MUX_SEL<='0';
																		 Rmadd<='0'&IR(8 DOWNTO 6);
																		 Rnadd<='0'&IR(5 DOWNTO 3);
																		 Rdadd<='0'&IR(2 DOWNTO 0);
																		 FLAGS<='1';
																		 CarryEn<='0';
																		 BIFURCATION<="0000";
																		 
													when "01110" => SEL<="00100";--ADD(immEDIATE)T1
																		 IMM<="00000000000000000000000000000"&IR(8 DOWNTO 6);
																		 MUX_SEL<='1';
																		 Rmadd<='0'&IR(5 DOWNTO 3);
																		 Rnadd<='0'&IR(5 DOWNTO 3);
																		 Rdadd<='0'&IR(2 DOWNTO 0);
																		 FLAGS<='1';
																		 CarryEn<='0';
																		 BIFURCATION<="0000";
																		 
													when "01111" => SEL<="00101";--SUB(immediate)T1
																		 IMM<="00000000000000000000000000000"&IR(8 DOWNTO 6);
																		 MUX_SEL<='1';
																		 Rmadd<='0'&IR(5 DOWNTO 3);
																		 Rnadd<='0'&IR(5 DOWNTO 3);
																		 Rdadd<='0'&IR(2 DOWNTO 0);
																		 FLAGS<='1';
																		 CarryEn<='0';
																		 BIFURCATION<="0000";
																		 
													when others => SEL<="ZZZZZ";
												END CASE;
														 
									when "100" => SEL<="10101";--MOV(immediate)
														 IMM<="000000000000000000000000"&IR(7 DOWNTO 0);
														 MUX_SEL<='1';
														 Rmadd<='0'&IR(5 DOWNTO 3);
														 Rnadd<='0'&IR(2 DOWNTO 0);
														 Rdadd<='0'&IR(10 DOWNTO 8);
														 FLAGS<='1';
														 CarryEn<='0';
														 BIFURCATION<="0000";
												
									when "101" => SEL<="00101";--CMP(immediate)
														 IMM<="000000000000000000000000"&IR(7 DOWNTO 0);
														 MUX_SEL<='1';
														 Rmadd<='0'&IR(10 DOWNTO 8);
														 Rnadd<='0'&IR(10 DOWNTO 8);
														 Rdadd<='0'&IR(2 DOWNTO 0);
														 FLAGS<='1';
														 CarryEn<='0';
														 BIFURCATION<="0001";
									
									when "110" => SEL<="00100";--ADD(immediate)T2
														 IMM<="000000000000000000000000"&IR(7 DOWNTO 0);
														 MUX_SEL<='1';
														 Rmadd<='0'&IR(10 DOWNTO 8);
														 Rnadd<='0'&IR(10 DOWNTO 8);
														 Rdadd<='0'&IR(10 DOWNTO 8);
														 FLAGS<='1';
														 CarryEn<='0';
														 BIFURCATION<="0000";
									
									when "111" => SEL<="00101";--SUB(immediate)T2
														 IMM<="000000000000000000000000"&IR(7 DOWNTO 0);
														 MUX_SEL<='1';
														 Rmadd<='0'&IR(5 DOWNTO 3);
														 Rnadd<='0'&IR(10 DOWNTO 8);
														 Rdadd<='0'&IR(10 DOWNTO 8);
														 FLAGS<='1';
														 CarryEn<='0';
														 BIFURCATION<="0000";
														 
									when others => SEL<="ZZZZZ"; 
								END CASE;
		
		when "01" =>
								CASE IR(13) IS
									WHEN '0' =>			
														CASE IR(12) IS
															WHEN '0' =>		
																			CASE IR(11 DOWNTO 10) IS
																				WHEN "00"=>
																								
																							 case IR(9 DOWNTO 6) is
																									when "0000" => SEL<="00000";--AND(register)
																														 MUX_SEL<='0';
																														 Rmadd<='0'&IR(5 DOWNTO 3);
																														 Rnadd<='0'&IR(2 DOWNTO 0);
																														 Rdadd<='0'&IR(2 DOWNTO 0);
																														 FLAGS<='1';
																														 CarryEn<='0';
																														 BIFURCATION<="0000";
																														 
																									when "0001" => SEL<="00010";--EOR(register)
																														 MUX_SEL<='0';
																														 Rmadd<='0'&IR(5 DOWNTO 3);
																														 Rnadd<='0'&IR(2 DOWNTO 0);
																														 Rdadd<='0'&IR(2 DOWNTO 0);
																														 FLAGS<='1';
																														 CarryEn<='0';
																														 BIFURCATION<="0000";
																									
																									when "0010" => SEL<="00110";--LSL(register)
																														 MUX_SEL<='0';
																														 Rmadd<='0'&IR(5 DOWNTO 3);
																														 Rnadd<='0'&IR(2 DOWNTO 0);
																														 Rdadd<='0'&IR(2 DOWNTO 0);
																														 FLAGS<='1';
																														 CarryEn<='0';
																														 BIFURCATION<="0000";
																									
																									when "0011" => SEL<="00111";--LSR(register)
																														 MUX_SEL<='0';
																														 Rmadd<='0'&IR(5 DOWNTO 3);
																														 Rnadd<='0'&IR(2 DOWNTO 0);
																														 Rdadd<='0'&IR(2 DOWNTO 0);
																														 FLAGS<='1';
																														 CarryEn<='0';
																														 BIFURCATION<="0000";
																									
																									when "0100" => SEL<="10000";--ASR(register)
																														 MUX_SEL<='0';
																														 Rmadd<='0'&IR(5 DOWNTO 3);
																														 Rnadd<='0'&IR(2 DOWNTO 0);
																														 Rdadd<='0'&IR(2 DOWNTO 0);
																														 FLAGS<='1';
																														 CarryEn<='0';
																														 BIFURCATION<="0000";
																														 
																									when "0101" => SEL<="00100";--ADC(register)
																														 MUX_SEL<='0';
																														 Rmadd<='0'&IR(5 DOWNTO 3);
																														 Rnadd<='0'&IR(2 DOWNTO 0);
																														 Rdadd<='0'&IR(2 DOWNTO 0);
																														 FLAGS<='1';
																														 CarryEn<='1';
																														 BIFURCATION<="0000";
																														 
																									when "0110" => SEL<="00101";--SBC(register)
																														 MUX_SEL<='0';
																														 Rmadd<='0'&IR(5 DOWNTO 3);
																														 Rnadd<='0'&IR(2 DOWNTO 0);
																														 Rdadd<='0'&IR(2 DOWNTO 0);
																														 FLAGS<='1';
																														 CarryEn<='1';
																														 BIFURCATION<="0000";
																														 
																									when "0111" => SEL<="10001";--ROR(register)
																														 MUX_SEL<='0';
																														 Rmadd<='0'&IR(5 DOWNTO 3);
																														 Rnadd<='0'&IR(2 DOWNTO 0);
																														 Rdadd<='0'&IR(2 DOWNTO 0);
																														 FLAGS<='1';
																														 CarryEn<='0';
																														 BIFURCATION<="0000";
																									
																									when "1000" => SEL<="00000";--TST(register)
																														 MUX_SEL<='0';
																														 Rmadd<='0'&IR(5 DOWNTO 3);
																														 Rnadd<='0'&IR(2 DOWNTO 0);
																														 Rdadd<='0'&IR(2 DOWNTO 0);
																														 FLAGS<='1';
																														 CarryEn<='0';
																														 BIFURCATION<="0001";
																									
																									when "1001" => SEL<="10110";--RSB(immediate)
																														 MUX_SEL<='0';
																														 Rmadd<='0'&IR(5 DOWNTO 3);
																														 Rnadd<='0'&IR(5 DOWNTO 3);
																														 Rdadd<='0'&IR(2 DOWNTO 0);
																														 FLAGS<='1';
																														 CarryEn<='0';
																														 BIFURCATION<="0000";
																									
																									when "1010" => SEL<="00101";--CMP(register)T1
																														 MUX_SEL<='0';
																														 Rmadd<='0'&IR(5 DOWNTO 3);
																														 Rnadd<='0'&IR(2 DOWNTO 0);
																														 Rdadd<='0'&IR(2 DOWNTO 0);
																														 FLAGS<='1';
																														 CarryEn<='0';
																														 BIFURCATION<="0001";
																									
																									when "1011" => SEL<="00100";--CMN(register)
																														 MUX_SEL<='0';
																														 Rmadd<='0'&IR(5 DOWNTO 3);
																														 Rnadd<='0'&IR(2 DOWNTO 0);
																														 Rdadd<='0'&IR(2 DOWNTO 0);
																														 FLAGS<='1';
																														 CarryEn<='0';
																														 BIFURCATION<="0001";
																														 
																									when "1100" => SEL<="00001";--ORR(register)
																														 MUX_SEL<='0';
																														 Rmadd<='0'&IR(5 DOWNTO 3);
																														 Rnadd<='0'&IR(2 DOWNTO 0);
																														 Rdadd<='0'&IR(2 DOWNTO 0);
																														 FLAGS<='1';
																														 CarryEn<='0';
																														 BIFURCATION<="0000";
																									
																									when "1101" => SEL<="10010";--MUL
																														 MUX_SEL<='0';
																														 Rmadd<='0'&IR(5 DOWNTO 3);
																														 Rnadd<='0'&IR(2 DOWNTO 0);
																														 Rdadd<='0'&IR(2 DOWNTO 0);
																														 FLAGS<='1';
																														 CarryEn<='0';
																														 BIFURCATION<="0010";
																									
																									when "1110" => SEL<="00011";--BIC(register)
																														 MUX_SEL<='0';
																														 Rmadd<='0'&IR(5 DOWNTO 3);
																														 Rnadd<='0'&IR(2 DOWNTO 0);
																														 Rdadd<='0'&IR(2 DOWNTO 0);
																														 FLAGS<='1';
																														 CarryEn<='0';
																														 BIFURCATION<="0000";
																														 
																									when "1111" => SEL<="10011";--MVN(register)
																														 MUX_SEL<='0';
																														 Rmadd<='0'&IR(5 DOWNTO 3);
																														 Rnadd<='0'&IR(5 DOWNTO 3);
																														 Rdadd<='0'&IR(2 DOWNTO 0);
																														 FLAGS<='1';
																														 CarryEn<='0';
																														 BIFURCATION<="0000";
																														 
																									WHEN OTHERS => SEL<="ZZZZZ";
																								END CASE;
																				
																				WHEN "01"=>	--Special data instructions and BRANCH and EXCHANGE		
																								
																								 case IR(9 DOWNTO 8) is
																									WHEN "00"=>
																													 SEL<="00100";--ADD(register)T2/ADD (SP PLUS REGISTER)T1/T2
																													 MUX_SEL<='0';
																													 Rmadd<=IR(6 DOWNTO 3);
																													 Rnadd<=IR(7)&IR(2 DOWNTO 0);
																													 Rdadd<=IR(7)&IR(2 DOWNTO 0);
																													 FLAGS<='0';
																													 CarryEn<='0';
																													 BIFURCATION<="0000";
																														 
																									WHEN "01"=>	SEL<="00101";--CMP(register)T2 
																													 MUX_SEL<='0';
																													 Rmadd<=IR(6 DOWNTO 3);
																													 Rnadd<=IR(7)&IR(2 DOWNTO 0);
																													 Rdadd<='1'&IR(2 DOWNTO 0);
																													 FLAGS<='1';
																													 CarryEn<='0';
																													 BIFURCATION<="0001";				
																													
																									WHEN "10"=>					
																													 SEL<="10101";--MOV(register)T1
																													 MUX_SEL<='0';
																													 Rmadd<=IR(6 DOWNTO 3);
																													 Rnadd<=IR(7)&IR(2 DOWNTO 0);
																													 Rdadd<=IR(7)&IR(2 DOWNTO 0);
																													 FLAGS<='0';
																													 CarryEn<='0';
																													 BIFURCATION<="0000";
																													 
																									WHEN "11"=>
																													CASE IR(7) IS	
																														when '0' => SEL<="10100";--BX 
																																			 MUX_SEL<='0';
																																			 Rmadd<=IR(6 DOWNTO 3);
																																			 Rnadd<=IR(6 DOWNTO 3);
																																			 Rdadd<="1111";
																																			 FLAGS<='0';
																																			 CarryEn<='0';
																																			 BIFURCATION<="0000";
																																			 
																														when '1' => --BLX(register)
																																			 
																																			 IMM<="00000000000000000000000000000001";
																																			 Rmadd<=IR(6 DOWNTO 3);
																																			 Rnadd<="1111";
																																			 FLAGS<='0';
																																			 CarryEn<='0';
																																			 BIFURCATION<="0110";
																																			 IF(FETCH1='1' OR FETCH2='1' OR FETCH3='1' OR BLX1='1' OR BLX2='1') THEN
																																					SEL<="00101";
																																					MUX_SEL<='1';
																																					Rdadd<="1110";
																																			  ELSE
																																					SEL<="10101";
																																					MUX_SEL<='0';
																																					Rdadd<="1111";
																																			  END IF;
																																			 
																														WHEN OTHERS=> SEL<="ZZZZZ";
																													END CASE;
																														
																									WHEN OTHERS=> SEL<="ZZZZZ";
																								END CASE;
																				WHEN "10"=>			
																							  SEL<="00100";--LDR(LITERAL)
																							  IMM<="000000000000000000000000"&IR(7 DOWNTO 0);
																							  MUX_SEL<='1';
																							  Rmadd<="1111";
																							  Rnadd<="1111";
																							  Rdadd<='0'&IR(10 DOWNTO 8);
																							  FLAGS<='0';
																							  CarryEn<='0';
																							  BIFURCATION<="0100";
																				
																				WHEN "11"=>			
																							  SEL<="00100";--LDR(LITERAL)
																							  IMM<="000000000000000000000000"&IR(7 DOWNTO 0);
																							  MUX_SEL<='1';
																							  Rmadd<="1111";
																							  Rnadd<="1111";
																							  Rdadd<='0'&IR(10 DOWNTO 8);
																							  FLAGS<='0';
																							  CarryEn<='0';
																							  BIFURCATION<="0100";
																							  
																				WHEN OTHERS => SEL<="ZZZZZ";
																			END CASE;
															WHEN '1'=>	--Load/store single data item				  
																				
																				 case IR(11 DOWNTO 9) is
																					when "000" => --STR(register) 
																										 MUX_SEL<='0';
																										 FLAGS<='0';
																										 CarryEn<='0';
																										 BIFURCATION<="0011";
																										 IF(FETCH1='1' OR FETCH2='1' OR FETCH3='1' OR STR1='1' OR STR2='1') THEN
																												SEL<="00100";
																												Rmadd<='0'&IR(8 DOWNTO 6);
																												Rnadd<='0'&IR(5 DOWNTO 3);
																												Rdadd<='0'&IR(2 DOWNTO 0);
																										  ELSE
																												SEL<="10100";
																												Rmadd<='0'&IR(2 DOWNTO 0);
																												Rnadd<='0'&IR(2 DOWNTO 0);
																												Rdadd<='0'&IR(2 DOWNTO 0);
																										  END IF;
																										 
																					
																					when "001" => --STRH(register) 
																										 MUX_SEL<='0';
																										 FLAGS<='0';
																										 CarryEn<='0';
																										 BIFURCATION<="0011";
																										 IF(FETCH1='1' OR FETCH2='1' OR FETCH3='1' OR STR1='1' OR STR2='1') THEN
																												SEL<="00100";
																												Rmadd<='0'&IR(8 DOWNTO 6);
																												Rnadd<='0'&IR(5 DOWNTO 3);
																												Rdadd<='0'&IR(2 DOWNTO 0);
																										  ELSE
																												SEL<="01010";
																												Rmadd<='0'&IR(2 DOWNTO 0);
																												Rnadd<='0'&IR(2 DOWNTO 0);
																												Rdadd<='0'&IR(2 DOWNTO 0);
																										  END IF;
																										 
																					when "010" => --STRB(register) 
																										 MUX_SEL<='0';
																										 FLAGS<='0';
																										 CarryEn<='0';
																										 BIFURCATION<="0011";
																										 IF(FETCH1='1' OR FETCH2='1' OR FETCH3='1' OR STR1='1' OR STR2='1') THEN
																												SEL<="00100";
																												Rmadd<='0'&IR(8 DOWNTO 6);
																												Rnadd<='0'&IR(5 DOWNTO 3);
																												Rdadd<='0'&IR(2 DOWNTO 0);
																										  ELSE
																												SEL<="01011";
																												Rmadd<='0'&IR(2 DOWNTO 0);
																												Rnadd<='0'&IR(2 DOWNTO 0);
																												Rdadd<='0'&IR(2 DOWNTO 0);
																										  END IF;
																										 
																					when "011" => --LDRSB(register)
																										 MUX_SEL<='0';
																										 FLAGS<='0';
																										 CarryEn<='0';
																										 BIFURCATION<="0101";
																										 IF(FETCH1='1' OR FETCH2='1' OR FETCH3='1' OR LOAD1='1' OR LOAD2='1') THEN
																												SEL<="00100";
																												Rmadd<='0'&IR(8 DOWNTO 6);
																												Rnadd<='0'&IR(5 DOWNTO 3);
																												Rdadd<='0'&IR(2 DOWNTO 0);
																										  ELSE
																												SEL<="01001";
																												Rmadd<='0'&IR(2 DOWNTO 0);
																												Rnadd<='0'&IR(2 DOWNTO 0);
																												Rdadd<='0'&IR(2 DOWNTO 0);
																										  END IF;
																							
																					when "100" => SEL<="00100";--LDR(register)
																										 MUX_SEL<='0';
																										 Rmadd<='0'&IR(8 DOWNTO 6);
																										 Rnadd<='0'&IR(5 DOWNTO 3);
																										 Rdadd<='0'&IR(2 DOWNTO 0);
																										 FLAGS<='0';
																										 CarryEn<='0';
																										 BIFURCATION<="0100";
																										 
																					when "101" => --LDRH(register) 
																										 MUX_SEL<='0';
																										 FLAGS<='0';
																										 CarryEn<='0';
																										 BIFURCATION<="0101";
																										 IF(FETCH1='1' OR FETCH2='1' OR FETCH3='1' OR LOAD1='1' OR LOAD2='1') THEN
																												SEL<="00100";
																												Rmadd<='0'&IR(8 DOWNTO 6);
																												Rnadd<='0'&IR(5 DOWNTO 3);
																												Rdadd<='0'&IR(2 DOWNTO 0);
																										  ELSE
																												SEL<="01010";
																												Rmadd<='0'&IR(2 DOWNTO 0);
																												Rnadd<='0'&IR(2 DOWNTO 0);
																												Rdadd<='0'&IR(2 DOWNTO 0);
																										  END IF;
																										 
																					when "110" => --LDRB(register)
																										 MUX_SEL<='0';
																										 FLAGS<='0';
																										 CarryEn<='0';
																										 BIFURCATION<="0101";
																										 IF(FETCH1='1' OR FETCH2='1' OR FETCH3='1' OR LOAD1='1' OR LOAD2='1') THEN
																												SEL<="00100";
																												Rmadd<='0'&IR(8 DOWNTO 6);
																												Rnadd<='0'&IR(5 DOWNTO 3);
																												Rdadd<='0'&IR(2 DOWNTO 0);
																										  ELSE
																												SEL<="01011";
																												Rmadd<='0'&IR(2 DOWNTO 0);
																												Rnadd<='0'&IR(2 DOWNTO 0);
																												Rdadd<='0'&IR(2 DOWNTO 0);
																										  END IF;
																					
																					when "111" => --LDRSH(register)
																										 MUX_SEL<='0';
																										 FLAGS<='0';
																										 CarryEn<='0';
																										 BIFURCATION<="0101";
																										 IF(FETCH1='1' OR FETCH2='1' OR FETCH3='1' OR LOAD1='1' OR LOAD2='1') THEN
																												SEL<="00100";
																												Rmadd<='0'&IR(8 DOWNTO 6);
																												Rnadd<='0'&IR(5 DOWNTO 3);
																												Rdadd<='0'&IR(2 DOWNTO 0);
																										  ELSE
																												SEL<="01000";
																												Rmadd<='0'&IR(2 DOWNTO 0);
																												Rnadd<='0'&IR(2 DOWNTO 0);
																												Rdadd<='0'&IR(2 DOWNTO 0);
																										  END IF;
																					
																					when others => SEL<="ZZZZZ";
																				END CASE;
															WHEN OTHERS=> SEL<="ZZZZZ";
														END CASE;
									WHEN '1' =>
															
														 case IR(12 DOWNTO 11) is
															when "00" => --STR(immediate)T1 
																				 IMM<="000000000000000000000000000"&IR(10 DOWNTO 6);
																				 MUX_SEL<='1';
																				 FLAGS<='0';
																				 CarryEn<='0';
																				 BIFURCATION<="0011";
																				 IF(FETCH1='1' OR FETCH2='1' OR FETCH3='1' OR STR1='1' OR STR2='1') THEN
																						SEL<="00100";
																						
																						Rmadd<='0'&IR(5 DOWNTO 3);
																						Rnadd<='0'&IR(5 DOWNTO 3);
																						Rdadd<='0'&IR(2 DOWNTO 0);
																				  ELSE
																						SEL<="10100";
																						--MUX_SEL<='0';
																						Rmadd<='0'&IR(2 DOWNTO 0);
																						Rnadd<='0'&IR(2 DOWNTO 0);
																						Rdadd<='0'&IR(2 DOWNTO 0);
																				  END IF;
															
															when "01" => SEL<="00100";--LDR(immEDIATE)T1 
																				 IMM<="000000000000000000000000000"&IR(10 DOWNTO 6);
																				 MUX_SEL<='1';
																				 Rmadd<='0'&IR(5 DOWNTO 3);
																				 Rnadd<='0'&IR(5 DOWNTO 3);
																				 Rdadd<='0'&IR(2 DOWNTO 0);
																				 FLAGS<='0';
																				 CarryEn<='0';
																				 BIFURCATION<="0100";
																				 
															when "10" => --STRB(IMMEDIATE) 
																				 IMM<="000000000000000000000000000"&IR(10 DOWNTO 6);
																				 FLAGS<='0';
																				 CarryEn<='0';
																				 BIFURCATION<="0011";
																				 IF(FETCH1='1' OR FETCH2='1' OR FETCH3='1' OR STR1='1' OR STR2='1') THEN
																						SEL<="00100";
																						MUX_SEL<='1';
																						Rmadd<='0'&IR(5 DOWNTO 3);
																						Rnadd<='0'&IR(5 DOWNTO 3);
																						Rdadd<='0'&IR(2 DOWNTO 0);
																				  ELSE
																						SEL<="01011";
																						MUX_SEL<='0';
																						Rmadd<='0'&IR(2 DOWNTO 0);
																						Rnadd<='0'&IR(2 DOWNTO 0);
																						Rdadd<='0'&IR(2 DOWNTO 0);
																				  END IF;
																				 
															when "11" => --LDRB(IMMEDIATE)
																				 IMM<="000000000000000000000000000"&IR(10 DOWNTO 6);
																				 FLAGS<='0';
																				 CarryEn<='0';
																				 BIFURCATION<="0101";
																				 IF(FETCH1='1' OR FETCH2='1' OR FETCH3='1' OR LOAD1='1' OR LOAD2='1') THEN
																						SEL<="00100";
																						MUX_SEL<='1';
																						Rmadd<='0'&IR(5 DOWNTO 3);
																						Rnadd<='0'&IR(5 DOWNTO 3);
																						Rdadd<='0'&IR(2 DOWNTO 0);
																				  ELSE
																						SEL<="01011";
																						MUX_SEL<='0';
																						Rmadd<='0'&IR(2 DOWNTO 0);
																						Rnadd<='0'&IR(2 DOWNTO 0);
																						Rdadd<='0'&IR(2 DOWNTO 0);
																				  END IF;
															
															WHEN OTHERS => SEL<="ZZZZZ";
														END CASE;
									WHEN OTHERS =>SEL<="ZZZZZ";
								END CASE; 
		WHEN "10"=>
						CASE IR(13) IS
							WHEN '0' =>--Load/store single data item
											 case IR(12 DOWNTO 11) is
												when "00" => --STRH(immediate) 
																	 IMM<="000000000000000000000000000"&IR(10 DOWNTO 6);
																	 FLAGS<='0';
																	 CarryEn<='0';
																	 BIFURCATION<="0011";
																	 IF(FETCH1='1' OR FETCH2='1' OR FETCH3='1' OR STR1='1' OR STR2='1') THEN
																			SEL<="00100";
																			MUX_SEL<='1';
																			Rmadd<='0'&IR(5 DOWNTO 3);
																			Rnadd<='0'&IR(5 DOWNTO 3);
																			Rdadd<='0'&IR(2 DOWNTO 0);
																	  ELSE
																			SEL<="01010";
																			MUX_SEL<='0';
																			Rmadd<='0'&IR(2 DOWNTO 0);
																			Rnadd<='0'&IR(2 DOWNTO 0);
																			Rdadd<='0'&IR(2 DOWNTO 0);
																	  END IF;
												
												when "01" => --LDRH(immEDIATE)
																	 IMM<="000000000000000000000000000"&IR(10 DOWNTO 6);
																	 FLAGS<='0';
																	 CarryEn<='0';
																	 BIFURCATION<="0101";
																	 IF(FETCH1='1' OR FETCH2='1' OR FETCH3='1' OR LOAD1='1' OR LOAD2='1') THEN
																			SEL<="00100";
																			MUX_SEL<='1';
																			Rmadd<='0'&IR(5 DOWNTO 3);
																			Rnadd<='0'&IR(5 DOWNTO 3);
																			Rdadd<='0'&IR(2 DOWNTO 0);
																	  ELSE
																			SEL<="01010";
																			MUX_SEL<='0';
																			Rmadd<='0'&IR(2 DOWNTO 0);
																			Rnadd<='0'&IR(2 DOWNTO 0);
																			Rdadd<='0'&IR(2 DOWNTO 0);
																	  END IF;
												
												when "10" => --STR(IMMEDIATE)T2 
																	 IMM<="000000000000000000000000"&IR(7 DOWNTO 0);
																	 FLAGS<='0';
																	 CarryEn<='0';
																	 BIFURCATION<="0011";
																	 IF(FETCH1='1' OR FETCH2='1' OR FETCH3='1' OR STR1='1' OR STR2='1') THEN
																			SEL<="00100";
																			MUX_SEL<='1';
																			Rmadd<="1101";
																			Rnadd<="1101";
																			Rdadd<="1101";
																	  ELSE
																			SEL<="10100";
																			MUX_SEL<='0';
																			Rmadd<='0'&IR(10 DOWNTO 8);
																			Rnadd<='0'&IR(10 DOWNTO 8);
																			Rdadd<='0'&IR(2 DOWNTO 0);
																	  END IF;
																	 
												when "11" => SEL<="00100";--LDR(IMMEDIATE)T2 
																	 IMM<="000000000000000000000000"&IR(7 DOWNTO 0);
																	 MUX_SEL<='1';
																	 Rmadd<="1101";
																	 Rnadd<="1101";
																	 Rdadd<='0'&IR(10 DOWNTO 8);
																	 FLAGS<='0';
																	 CarryEn<='0';
																	 BIFURCATION<="0100";
												
												WHEN OTHERS => SEL<="ZZZZZ";
											END CASE;
							WHEN '1'=>
											CASE IR(12) IS
												WHEN '0'=>
																CASE IR(11) IS
																	WHEN '0'=>
																				  SEL<="00100";--ADR
																				  IMM<="000000000000000000000000"&IR(7 DOWNTO 0);
																				  MUX_SEL<='1';
																				  Rmadd<="1111";
																				  Rnadd<="1111";
																				  Rdadd<='0'&IR(10 DOWNTO 8);
																				  FLAGS<='0';
																				  CarryEn<='0';
																				  BIFURCATION<="0000";
																				  
																	WHEN '1'=>		
																				  SEL<="00100";--ADD(SP PLUS IMMEDIATE)T1
																				  IMM<="000000000000000000000000"&IR(7 DOWNTO 0);
																				  MUX_SEL<='1';
																				  Rmadd<="1101";
																				  Rnadd<="1101";
																				  Rdadd<='0'&IR(10 DOWNTO 8);
																				  FLAGS<='0';
																				  CarryEn<='0';
																				  BIFURCATION<="0000";
																				  
																	WHEN OTHERS=>SEL<="ZZZZZ";
																END CASE;
												
												WHEN '1'=>--Load/store single data item		
																
																 case IR(11 DOWNTO 9) is
																	WHEN "000"=>	
																						case IR(11 DOWNTO 7) is
																							when "00000" => SEL<="00100";--ADD(SP PLUS IMMEDIATE)T2
																												 IMM<="0000000000000000000000000"&IR(6 DOWNTO 0);
																												 MUX_SEL<='1';
																												 Rmadd<="1101";
																												 Rnadd<="1101";
																												 Rdadd<="1101";
																												 FLAGS<='0';
																												 CarryEn<='0';
																												 BIFURCATION<="0000";
																							
																							when "00001" => SEL<="00101";--SUB(SP minus IMMEDIATE)T1 
																												 IMM<="0000000000000000000000000"&IR(6 DOWNTO 0);
																												 MUX_SEL<='1';
																												 Rmadd<=IR(6 DOWNTO 3);
																												 Rnadd<="1101";
																												 Rdadd<="1101";
																												 FLAGS<='0';
																												 CarryEn<='0';
																												 BIFURCATION<="0000";
																												 
																							WHEN OTHERS => SEL<="ZZZZZ";
																						END CASE;
																	WHEN "001"=>					
																					case IR(11 DOWNTO 6) is
																						when "001000" => SEL<="01000";--SXTH
																											 MUX_SEL<='0';
																											 Rmadd<='0'&IR(5 DOWNTO 3);
																											 Rnadd<='0'&IR(5 DOWNTO 3);
																											 Rdadd<='0'&IR(2 DOWNTO 0);
																											 FLAGS<='0';
																											 CarryEn<='0';
																											 BIFURCATION<="0000";
																											 
																						when "001001" => SEL<="01001";--SXTB 
																											 MUX_SEL<='0';
																											 Rmadd<='0'&IR(5 DOWNTO 3);
																											 Rnadd<='0'&IR(5 DOWNTO 3);
																											 Rdadd<='0'&IR(2 DOWNTO 0);
																											 FLAGS<='0';
																											 CarryEn<='0';
																											 BIFURCATION<="0000";
																						
																						when "001010" => SEL<="01010";--UXTH
																											 MUX_SEL<='0';
																											 Rmadd<='0'&IR(5 DOWNTO 3);
																											 Rnadd<='0'&IR(5 DOWNTO 3);
																											 Rdadd<='0'&IR(2 DOWNTO 0);
																											 FLAGS<='0';
																											 CarryEn<='0';
																											 BIFURCATION<="0000";
																											 
																						when "001011" => SEL<="01011";--UXTB 
																											 MUX_SEL<='0';
																											 Rmadd<='0'&IR(5 DOWNTO 3);
																											 Rnadd<='0'&IR(5 DOWNTO 3);
																											 Rdadd<='0'&IR(2 DOWNTO 0);
																											 FLAGS<='0';
																											 CarryEn<='0';
																											 BIFURCATION<="0000";
																											 
																						WHEN OTHERS=> SEL<="ZZZZZ";
																					END CASE;
																					
																	WHEN "010"=>--PUSH 
																				 IMM<="00000000000000000000000000000100";
																				 MUX_SEL<='1';
																				 FLAGS<='0';
																				 CarryEn<='0';
																				 BIFURCATION<="1000";
																				 IF(FETCH1='1' OR FETCH2='1' OR FETCH3='1' OR PUSH1='1' OR PUSH2='1'OR PUSH6='1' OR PUSH7='1' OR
																					 PUSH11='1' OR PUSH12='1' OR PUSH16='1' OR PUSH17='1' OR PUSH21='1' OR PUSH22='1' OR
																					 PUSH26='1' OR PUSH27='1' OR PUSH31='1' OR PUSH32='1' OR PUSH36='1' OR PUSH37='1' OR
																					 PUSH41='1' OR PUSH42='1') THEN
																						SEL<="00100";
																					   Rmadd<="1110";
																						Rnadd<="1110";
																						Rdadd<="1110";
																				  ELSIF(PUSH3='1' OR PUSH4='1' OR PUSH5='1')THEN 
																						SEL<="10100";
																						Rmadd<="0000";
																						Rnadd<="0000";
																						Rdadd<="0000";
																				  ELSIF(PUSH8='1' OR PUSH9='1' OR PUSH10='1')THEN 
																						SEL<="10100";
																						Rmadd<="0001";
																						Rnadd<="0001";
																						Rdadd<="0001";
																				  ELSIF(PUSH13='1' OR PUSH14='1' OR PUSH15='1')THEN 
																						SEL<="10100";
																						Rmadd<="0010";
																						Rnadd<="0010";
																						Rdadd<="0010";
																				  ELSIF(PUSH18='1' OR PUSH19='1' OR PUSH20='1')THEN 
																						SEL<="10100";
																						Rmadd<="0011";
																						Rnadd<="0011";
																						Rdadd<="0011";
																				  ELSIF(PUSH23='1' OR PUSH24='1' OR PUSH25='1')THEN 
																						SEL<="10100";
																						Rmadd<="0100";
																						Rnadd<="0100";
																						Rdadd<="0100";
																				  ELSIF(PUSH28='1' OR PUSH29='1' OR PUSH30='1')THEN 
																						SEL<="10100";
																						Rmadd<="0101";
																						Rnadd<="0101";
																						Rdadd<="0101";
																				  ELSIF(PUSH33='1' OR PUSH34='1' OR PUSH35='1')THEN 
																						SEL<="10100";
																						Rmadd<="0110";
																						Rnadd<="0110";
																						Rdadd<="0110";
																				  ELSIF(PUSH38='1' OR PUSH39='1' OR PUSH40='1')THEN 
																						SEL<="10100";
																						Rmadd<="0111";
																						Rnadd<="0111";
																						Rdadd<="0111";
																				  ELSIF(PUSH43='1' OR PUSH44='1' OR PUSH45='1')THEN 
																						SEL<="10100";
																						Rmadd<="1101";
																						Rnadd<="1101";
																						Rdadd<="1101";
																					ELSE NULL;
																				  END IF;
																					 
																					 
																	WHEN "101"=>										 
																					CASE IR(11 DOWNTO 6) IS	
																						when "101000" => SEL<="01100";--REV 
																											 MUX_SEL<='0';
																											 Rmadd<='0'&IR(5 DOWNTO 3);
																											 Rnadd<='0'&IR(5 DOWNTO 3);
																											 Rdadd<='0'&IR(2 DOWNTO 0);
																											 FLAGS<='0';
																											 CarryEn<='0';
																											 BIFURCATION<="0000";
																						
																						when "101001" => SEL<="01101";--REV16
																											 MUX_SEL<='0';
																											 Rmadd<='0'&IR(5 DOWNTO 3);
																											 Rnadd<='0'&IR(5 DOWNTO 3);
																											 Rdadd<='0'&IR(2 DOWNTO 0);
																											 FLAGS<='0';
																											 CarryEn<='0';
																											 BIFURCATION<="0000";
																											 
																						when "101011" => SEL<="01111";--REVSH 
																											 MUX_SEL<='0';
																											 Rmadd<='0'&IR(5 DOWNTO 3);
																											 Rnadd<='0'&IR(5 DOWNTO 3);
																											 Rdadd<='0'&IR(2 DOWNTO 0);
																											 FLAGS<='0';
																											 CarryEn<='0';
																											 BIFURCATION<="0000";
																											 
																						WHEN OTHERS=> SEL<="ZZZZZ";
																					END CASE;
																	WHEN "110"=>--POP 
																				 IMM<="00000000000000000000000000000100"; 
																				 MUX_SEL<='1';
																				 FLAGS<='0';
																				 CarryEn<='0';
																				 BIFURCATION<="1001";
																				 IF(FETCH1='1' OR FETCH2='1' OR FETCH3='1' OR POP1='1' OR POP2='1'  ) THEN
																						
																						SEL<="00100";
																					   Rmadd<="1110";
																						Rnadd<="1110";
																						Rdadd<="1110";
																				  ELSIF(POP3='1' OR POP4='1' OR POP7='1' OR POP8='1'OR POP11='1' OR POP12='1' OR
																					 POP15='1' OR POP16='1' OR POP19='1' OR POP20='1' OR POP23='1' OR POP24='1' OR
																					 POP27='1' OR POP28='1' OR POP31='1' OR POP32='1' OR POP35='1' OR POP36='1')THEN 
																						SEL<="00101";
																					   Rmadd<="1110";
																						Rnadd<="1110";
																						Rdadd<="1110";
																				  ELSIF(POP5='1' OR POP6='1')THEN 
																						SEL<="10100";
																						Rmadd<="0000";
																						Rnadd<="0000";
																						Rdadd<="0000";
																				  ELSIF(POP9='1' OR POP10='1')THEN 
																						SEL<="10100";
																						Rmadd<="0001";
																						Rnadd<="0001";
																						Rdadd<="0001";
																				  ELSIF(POP13='1' OR POP14='1')THEN 
																						SEL<="10100";
																						Rmadd<="0010";
																						Rnadd<="0010";
																						Rdadd<="0010";
																				  ELSIF(POP17='1' OR POP18='1')THEN 
																						SEL<="10100";
																						Rmadd<="0011";
																						Rnadd<="0011";
																						Rdadd<="0011";
																				  ELSIF(POP21='1' OR POP22='1')THEN 
																						SEL<="10100";
																						Rmadd<="0100";
																						Rnadd<="0100";
																						Rdadd<="0100";
																				  ELSIF(POP25='1' OR POP26='1')THEN 
																						SEL<="10100";
																						Rmadd<="0101";
																						Rnadd<="0101";
																						Rdadd<="0101";
																				  ELSIF(POP29='1' OR POP30='1')THEN 
																						SEL<="10100";
																						Rmadd<="0110";
																						Rnadd<="0110";
																						Rdadd<="0110";
																				  ELSIF(POP33='1' OR POP34='1')THEN 
																						SEL<="10100";
																						Rmadd<="0111";
																						Rnadd<="0111";
																						Rdadd<="0111";
																				  ELSIF(POP37='1' OR POP38='1')THEN 
																						SEL<="10100";
																						Rmadd<="1101";
																						Rnadd<="1101";
																						Rdadd<="1101";
																					ELSE NULL;
																				  END IF;
																	
																	WHEN "111"=>										 
																					 SEL<="11111";--NOP
																					 MUX_SEL<='0';
																					 Rmadd<='0'&IR(5 DOWNTO 3);
																					 Rnadd<='0'&IR(5 DOWNTO 3);
																					 Rdadd<='0'&IR(2 DOWNTO 0);
																					 FLAGS<='0';
																					 CarryEn<='0';
																					 BIFURCATION<="0001";
														
																	WHEN OTHERS => SEL<="ZZZZZ";
																END CASE;
												WHEN OTHERS=> SEL<="ZZZZZ";
											END CASE;
											
							WHEN OTHERS=> SEL<="ZZZZZ";
						END CASE;
		
		WHEN "11"=>
					CASE IR(13 DOWNTO 12) IS	
						when "01" => SEL<="00100";--B T1 
											 IMM<="000000000000000000000000"&IR(7 DOWNTO 0);
											 MUX_SEL<='1';
											 Rmadd<="1111";
											 Rnadd<="1111";
											 Rdadd<="1111";
											 FLAGS<='0';
											 CarryEn<='0';
											BIFURCATION<="0000";
											
--											IF ((IR(11 DOWNTO 8)="0000" AND NZCV(2)='1') OR 
--												 (IR(11 DOWNTO 8)="0001" AND NZCV(2)='0') OR
--												 (IR(11 DOWNTO 8)="0010" AND NZCV(1)='1') OR
--												 (IR(11 DOWNTO 8)="0011" AND NZCV(1)='0') OR
--												 (IR(11 DOWNTO 8)="0100" AND NZCV(3)='1') OR
--												 (IR(11 DOWNTO 8)="0101" AND NZCV(3)='0') OR
--												 (IR(11 DOWNTO 8)="0110" AND NZCV(0)='1') OR
--												 (IR(11 DOWNTO 8)="0111" AND NZCV(0)='0') OR
--												 (IR(11 DOWNTO 8)="1000" AND NZCV(1)='1' AND NZCV(2)='0') OR
--												 (IR(11 DOWNTO 8)="1001" AND (NZCV(1)='0' OR NZCV(2)='1')) OR
--												 (IR(11 DOWNTO 8)="1010" AND NZCV(3)=NZCV(0)) OR
--												 (IR(11 DOWNTO 8)="1011" AND ((NZCV(3)='1' AND NZCV(0)='0') OR (NZCV(3)='0' AND NZCV(0)='1'))) OR
--												 (IR(11 DOWNTO 8)="1100" AND NZCV(2)='0' AND NZCV(3)=NZCV(0)) OR
--												 (IR(11 DOWNTO 8)="1101" AND (NZCV(2)='1' OR (NZCV(3)='1' AND NZCV(0)='0') OR (NZCV(3)='0' AND NZCV(0)='1'))) OR
--												 IR(11 DOWNTO 8)="1110" OR IR(11 DOWNTO 8)="1111"
--											)THEN
--												BIFURCATION<="0000";
--											ELSE
--												BIFURCATION<="0001";
--											END IF;
											
					
									
											 
						when "10" => SEL<="00100";--B T2
											 MUX_SEL<='1';
											 IMM<="000000000000000000000"&IR(10 DOWNTO 0);
											 Rmadd<="1111";
											 Rnadd<="1111";
											 Rdadd<="1111";
											 FLAGS<='0';
											 CarryEn<='0';
											 BIFURCATION<="0000";
						
						when "11" => --BL 
											 
											 Rmadd<="1111";
											 Rnadd<="1111";
											 FLAGS<='0';
											 CarryEn<='0';
											 BIFURCATION<="0111";
											 IF(FETCH1='1' OR FETCH2='1' OR FETCH3='1' OR BL1='1' OR BL2='1') THEN
													MUX_SEL<='0';
													SEL<="10100";
													Rdadd<="1110";
											  ELSE
													MUX_SEL<='1';
													IMM<="0000000"&IR(10)&(IR(10) XOR IR2(13))&(IR(10)XOR IR2(11))&IR(9 DOWNTO 0)&IR2(10 DOWNTO 0)&'0';
													SEL<="10101";
													Rdadd<="1111";
											  END IF;
											 
						WHEN OTHERS=> SEL<="ZZZZZ";
						END CASE;
			
		WHEN OTHERS =>SEL<="ZZZZZ";
	END CASE;

END PROCESS;





end RTL;